[translated]
module main

pub struct Rectangle {
pub mut:
height any
length any
}

fn (self Rectangle) __init__ (height A, length B) {
    self.height = height
    self.length = length
}
fn main () {
    r := Rectangle{}
}
