[translated]
module main

{1: 1}.keys()
