[translated]
module main

pub struct A {

}

B := "FOO"
fn main () {
    assert A.B == "FOO"
}
